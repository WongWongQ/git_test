﻿module fpga(
		input		clk,
		input		rst_n,
		output a
		);
		
	endmodule